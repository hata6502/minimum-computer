module character_rom (
    input wire clock,
    input wire [2:0] x,
    input wire [2:0] y,
    input wire [6:0] character,
    output wire dot
);
  reg [7:0] character_line_data;

  assign dot = character_line_data[7-x];

  initial begin
    character_line_data = 0;
  end

  always @(posedge clock) begin
    case ({
      character, y
    })
      0: character_line_data <= 'b00000000;
      1: character_line_data <= 'b00000000;
      2: character_line_data <= 'b00000000;
      3: character_line_data <= 'b00000000;
      4: character_line_data <= 'b00000000;
      5: character_line_data <= 'b00000000;
      6: character_line_data <= 'b00000000;
      7: character_line_data <= 'b00000000;
      8: character_line_data <= 'b00000000;
      9: character_line_data <= 'b00000000;
      10: character_line_data <= 'b00000000;
      11: character_line_data <= 'b00000000;
      12: character_line_data <= 'b00000000;
      13: character_line_data <= 'b00000000;
      14: character_line_data <= 'b00000000;
      15: character_line_data <= 'b00000000;
      16: character_line_data <= 'b00000000;
      17: character_line_data <= 'b00000000;
      18: character_line_data <= 'b00000000;
      19: character_line_data <= 'b00000000;
      20: character_line_data <= 'b00000000;
      21: character_line_data <= 'b00000000;
      22: character_line_data <= 'b00000000;
      23: character_line_data <= 'b00000000;
      24: character_line_data <= 'b00000000;
      25: character_line_data <= 'b00000000;
      26: character_line_data <= 'b00000000;
      27: character_line_data <= 'b00000000;
      28: character_line_data <= 'b00000000;
      29: character_line_data <= 'b00000000;
      30: character_line_data <= 'b00000000;
      31: character_line_data <= 'b00000000;
      32: character_line_data <= 'b00000000;
      33: character_line_data <= 'b00000000;
      34: character_line_data <= 'b00000000;
      35: character_line_data <= 'b00000000;
      36: character_line_data <= 'b00000000;
      37: character_line_data <= 'b00000000;
      38: character_line_data <= 'b00000000;
      39: character_line_data <= 'b00000000;
      40: character_line_data <= 'b00000000;
      41: character_line_data <= 'b00000000;
      42: character_line_data <= 'b00000000;
      43: character_line_data <= 'b00000000;
      44: character_line_data <= 'b00000000;
      45: character_line_data <= 'b00000000;
      46: character_line_data <= 'b00000000;
      47: character_line_data <= 'b00000000;
      48: character_line_data <= 'b00000000;
      49: character_line_data <= 'b00000000;
      50: character_line_data <= 'b00000000;
      51: character_line_data <= 'b00000000;
      52: character_line_data <= 'b00000000;
      53: character_line_data <= 'b00000000;
      54: character_line_data <= 'b00000000;
      55: character_line_data <= 'b00000000;
      56: character_line_data <= 'b00000000;
      57: character_line_data <= 'b00000000;
      58: character_line_data <= 'b00000000;
      59: character_line_data <= 'b00000000;
      60: character_line_data <= 'b00000000;
      61: character_line_data <= 'b00000000;
      62: character_line_data <= 'b00000000;
      63: character_line_data <= 'b00000000;
      64: character_line_data <= 'b00000000;
      65: character_line_data <= 'b00000000;
      66: character_line_data <= 'b00000000;
      67: character_line_data <= 'b00000000;
      68: character_line_data <= 'b00000000;
      69: character_line_data <= 'b00000000;
      70: character_line_data <= 'b00000000;
      71: character_line_data <= 'b00000000;
      72: character_line_data <= 'b00000000;
      73: character_line_data <= 'b00000000;
      74: character_line_data <= 'b00000000;
      75: character_line_data <= 'b00000000;
      76: character_line_data <= 'b00000000;
      77: character_line_data <= 'b00000000;
      78: character_line_data <= 'b00000000;
      79: character_line_data <= 'b00000000;
      80: character_line_data <= 'b00000000;
      81: character_line_data <= 'b00000000;
      82: character_line_data <= 'b00000000;
      83: character_line_data <= 'b00000000;
      84: character_line_data <= 'b00000000;
      85: character_line_data <= 'b00000000;
      86: character_line_data <= 'b00000000;
      87: character_line_data <= 'b00000000;
      88: character_line_data <= 'b00000000;
      89: character_line_data <= 'b00000000;
      90: character_line_data <= 'b00000000;
      91: character_line_data <= 'b00000000;
      92: character_line_data <= 'b00000000;
      93: character_line_data <= 'b00000000;
      94: character_line_data <= 'b00000000;
      95: character_line_data <= 'b00000000;
      96: character_line_data <= 'b00000000;
      97: character_line_data <= 'b00000000;
      98: character_line_data <= 'b00000000;
      99: character_line_data <= 'b00000000;
      100: character_line_data <= 'b00000000;
      101: character_line_data <= 'b00000000;
      102: character_line_data <= 'b00000000;
      103: character_line_data <= 'b00000000;
      104: character_line_data <= 'b00000000;
      105: character_line_data <= 'b00000000;
      106: character_line_data <= 'b00000000;
      107: character_line_data <= 'b00000000;
      108: character_line_data <= 'b00000000;
      109: character_line_data <= 'b00000000;
      110: character_line_data <= 'b00000000;
      111: character_line_data <= 'b00000000;
      112: character_line_data <= 'b00000000;
      113: character_line_data <= 'b00000000;
      114: character_line_data <= 'b00000000;
      115: character_line_data <= 'b00000000;
      116: character_line_data <= 'b00000000;
      117: character_line_data <= 'b00000000;
      118: character_line_data <= 'b00000000;
      119: character_line_data <= 'b00000000;
      120: character_line_data <= 'b00000000;
      121: character_line_data <= 'b00000000;
      122: character_line_data <= 'b00000000;
      123: character_line_data <= 'b00000000;
      124: character_line_data <= 'b00000000;
      125: character_line_data <= 'b00000000;
      126: character_line_data <= 'b00000000;
      127: character_line_data <= 'b00000000;
      128: character_line_data <= 'b00000000;
      129: character_line_data <= 'b00000000;
      130: character_line_data <= 'b00000000;
      131: character_line_data <= 'b00000000;
      132: character_line_data <= 'b00000000;
      133: character_line_data <= 'b00000000;
      134: character_line_data <= 'b00000000;
      135: character_line_data <= 'b00000000;
      136: character_line_data <= 'b00000000;
      137: character_line_data <= 'b00000000;
      138: character_line_data <= 'b00000000;
      139: character_line_data <= 'b00000000;
      140: character_line_data <= 'b00000000;
      141: character_line_data <= 'b00000000;
      142: character_line_data <= 'b00000000;
      143: character_line_data <= 'b00000000;
      144: character_line_data <= 'b00000000;
      145: character_line_data <= 'b00000000;
      146: character_line_data <= 'b00000000;
      147: character_line_data <= 'b00000000;
      148: character_line_data <= 'b00000000;
      149: character_line_data <= 'b00000000;
      150: character_line_data <= 'b00000000;
      151: character_line_data <= 'b00000000;
      152: character_line_data <= 'b00000000;
      153: character_line_data <= 'b00000000;
      154: character_line_data <= 'b00000000;
      155: character_line_data <= 'b00000000;
      156: character_line_data <= 'b00000000;
      157: character_line_data <= 'b00000000;
      158: character_line_data <= 'b00000000;
      159: character_line_data <= 'b00000000;
      160: character_line_data <= 'b00000000;
      161: character_line_data <= 'b00000000;
      162: character_line_data <= 'b00000000;
      163: character_line_data <= 'b00000000;
      164: character_line_data <= 'b00000000;
      165: character_line_data <= 'b00000000;
      166: character_line_data <= 'b00000000;
      167: character_line_data <= 'b00000000;
      168: character_line_data <= 'b00000000;
      169: character_line_data <= 'b00000000;
      170: character_line_data <= 'b00000000;
      171: character_line_data <= 'b00000000;
      172: character_line_data <= 'b00000000;
      173: character_line_data <= 'b00000000;
      174: character_line_data <= 'b00000000;
      175: character_line_data <= 'b00000000;
      176: character_line_data <= 'b00000000;
      177: character_line_data <= 'b00000000;
      178: character_line_data <= 'b00000000;
      179: character_line_data <= 'b00000000;
      180: character_line_data <= 'b00000000;
      181: character_line_data <= 'b00000000;
      182: character_line_data <= 'b00000000;
      183: character_line_data <= 'b00000000;
      184: character_line_data <= 'b00000000;
      185: character_line_data <= 'b00000000;
      186: character_line_data <= 'b00000000;
      187: character_line_data <= 'b00000000;
      188: character_line_data <= 'b00000000;
      189: character_line_data <= 'b00000000;
      190: character_line_data <= 'b00000000;
      191: character_line_data <= 'b00000000;
      192: character_line_data <= 'b00000000;
      193: character_line_data <= 'b00000000;
      194: character_line_data <= 'b00000000;
      195: character_line_data <= 'b00000000;
      196: character_line_data <= 'b00000000;
      197: character_line_data <= 'b00000000;
      198: character_line_data <= 'b00000000;
      199: character_line_data <= 'b00000000;
      200: character_line_data <= 'b00000000;
      201: character_line_data <= 'b00000000;
      202: character_line_data <= 'b00000000;
      203: character_line_data <= 'b00000000;
      204: character_line_data <= 'b00000000;
      205: character_line_data <= 'b00000000;
      206: character_line_data <= 'b00000000;
      207: character_line_data <= 'b00000000;
      208: character_line_data <= 'b00000000;
      209: character_line_data <= 'b00000000;
      210: character_line_data <= 'b00000000;
      211: character_line_data <= 'b00000000;
      212: character_line_data <= 'b00000000;
      213: character_line_data <= 'b00000000;
      214: character_line_data <= 'b00000000;
      215: character_line_data <= 'b00000000;
      216: character_line_data <= 'b00000000;
      217: character_line_data <= 'b00000000;
      218: character_line_data <= 'b00000000;
      219: character_line_data <= 'b00000000;
      220: character_line_data <= 'b00000000;
      221: character_line_data <= 'b00000000;
      222: character_line_data <= 'b00000000;
      223: character_line_data <= 'b00000000;
      224: character_line_data <= 'b00000000;
      225: character_line_data <= 'b00000000;
      226: character_line_data <= 'b00000000;
      227: character_line_data <= 'b00000000;
      228: character_line_data <= 'b00000000;
      229: character_line_data <= 'b00000000;
      230: character_line_data <= 'b00000000;
      231: character_line_data <= 'b00000000;
      232: character_line_data <= 'b00000000;
      233: character_line_data <= 'b00000000;
      234: character_line_data <= 'b00000000;
      235: character_line_data <= 'b00000000;
      236: character_line_data <= 'b00000000;
      237: character_line_data <= 'b00000000;
      238: character_line_data <= 'b00000000;
      239: character_line_data <= 'b00000000;
      240: character_line_data <= 'b00000000;
      241: character_line_data <= 'b00000000;
      242: character_line_data <= 'b00000000;
      243: character_line_data <= 'b00000000;
      244: character_line_data <= 'b00000000;
      245: character_line_data <= 'b00000000;
      246: character_line_data <= 'b00000000;
      247: character_line_data <= 'b00000000;
      248: character_line_data <= 'b00000000;
      249: character_line_data <= 'b00000000;
      250: character_line_data <= 'b00000000;
      251: character_line_data <= 'b00000000;
      252: character_line_data <= 'b00000000;
      253: character_line_data <= 'b00000000;
      254: character_line_data <= 'b00000000;
      255: character_line_data <= 'b00000000;
      256: character_line_data <= 'b00000000;
      257: character_line_data <= 'b00000000;
      258: character_line_data <= 'b00000000;
      259: character_line_data <= 'b00000000;
      260: character_line_data <= 'b00000000;
      261: character_line_data <= 'b00000000;
      262: character_line_data <= 'b00000000;
      263: character_line_data <= 'b00000000;
      264: character_line_data <= 'b00010000;
      265: character_line_data <= 'b00010000;
      266: character_line_data <= 'b00010000;
      267: character_line_data <= 'b00010000;
      268: character_line_data <= 'b00010000;
      269: character_line_data <= 'b00000000;
      270: character_line_data <= 'b00010000;
      271: character_line_data <= 'b00000000;
      272: character_line_data <= 'b11011000;
      273: character_line_data <= 'b01001000;
      274: character_line_data <= 'b10010000;
      275: character_line_data <= 'b00000000;
      276: character_line_data <= 'b00000000;
      277: character_line_data <= 'b00000000;
      278: character_line_data <= 'b00000000;
      279: character_line_data <= 'b00000000;
      280: character_line_data <= 'b00010100;
      281: character_line_data <= 'b01111110;
      282: character_line_data <= 'b00101000;
      283: character_line_data <= 'b00101000;
      284: character_line_data <= 'b00101000;
      285: character_line_data <= 'b11111100;
      286: character_line_data <= 'b01010000;
      287: character_line_data <= 'b00000000;
      288: character_line_data <= 'b00001000;
      289: character_line_data <= 'b00111110;
      290: character_line_data <= 'b01001000;
      291: character_line_data <= 'b00111100;
      292: character_line_data <= 'b00010010;
      293: character_line_data <= 'b01111100;
      294: character_line_data <= 'b00010000;
      295: character_line_data <= 'b00000000;
      296: character_line_data <= 'b01000010;
      297: character_line_data <= 'b10100100;
      298: character_line_data <= 'b01001000;
      299: character_line_data <= 'b00010000;
      300: character_line_data <= 'b00100100;
      301: character_line_data <= 'b01001010;
      302: character_line_data <= 'b10000100;
      303: character_line_data <= 'b00000000;
      304: character_line_data <= 'b00110000;
      305: character_line_data <= 'b01001000;
      306: character_line_data <= 'b01010000;
      307: character_line_data <= 'b00100100;
      308: character_line_data <= 'b01010100;
      309: character_line_data <= 'b10001000;
      310: character_line_data <= 'b01110110;
      311: character_line_data <= 'b00000000;
      312: character_line_data <= 'b11000000;
      313: character_line_data <= 'b01000000;
      314: character_line_data <= 'b10000000;
      315: character_line_data <= 'b00000000;
      316: character_line_data <= 'b00000000;
      317: character_line_data <= 'b00000000;
      318: character_line_data <= 'b00000000;
      319: character_line_data <= 'b00000000;
      320: character_line_data <= 'b00000010;
      321: character_line_data <= 'b00000100;
      322: character_line_data <= 'b00001000;
      323: character_line_data <= 'b00001000;
      324: character_line_data <= 'b00001000;
      325: character_line_data <= 'b00000100;
      326: character_line_data <= 'b00000010;
      327: character_line_data <= 'b00000000;
      328: character_line_data <= 'b10000000;
      329: character_line_data <= 'b01000000;
      330: character_line_data <= 'b00100000;
      331: character_line_data <= 'b00100000;
      332: character_line_data <= 'b00100000;
      333: character_line_data <= 'b01000000;
      334: character_line_data <= 'b10000000;
      335: character_line_data <= 'b00000000;
      336: character_line_data <= 'b00010000;
      337: character_line_data <= 'b01010100;
      338: character_line_data <= 'b00111000;
      339: character_line_data <= 'b00010000;
      340: character_line_data <= 'b00111000;
      341: character_line_data <= 'b01010100;
      342: character_line_data <= 'b00010000;
      343: character_line_data <= 'b00000000;
      344: character_line_data <= 'b00010000;
      345: character_line_data <= 'b00010000;
      346: character_line_data <= 'b00010000;
      347: character_line_data <= 'b11111110;
      348: character_line_data <= 'b00010000;
      349: character_line_data <= 'b00010000;
      350: character_line_data <= 'b00010000;
      351: character_line_data <= 'b00000000;
      352: character_line_data <= 'b00000000;
      353: character_line_data <= 'b00000000;
      354: character_line_data <= 'b00000000;
      355: character_line_data <= 'b00000000;
      356: character_line_data <= 'b11000000;
      357: character_line_data <= 'b01000000;
      358: character_line_data <= 'b10000000;
      359: character_line_data <= 'b00000000;
      360: character_line_data <= 'b00000000;
      361: character_line_data <= 'b00000000;
      362: character_line_data <= 'b00000000;
      363: character_line_data <= 'b11111110;
      364: character_line_data <= 'b00000000;
      365: character_line_data <= 'b00000000;
      366: character_line_data <= 'b00000000;
      367: character_line_data <= 'b00000000;
      368: character_line_data <= 'b00000000;
      369: character_line_data <= 'b00000000;
      370: character_line_data <= 'b00000000;
      371: character_line_data <= 'b00000000;
      372: character_line_data <= 'b00000000;
      373: character_line_data <= 'b11000000;
      374: character_line_data <= 'b11000000;
      375: character_line_data <= 'b00000000;
      376: character_line_data <= 'b00000010;
      377: character_line_data <= 'b00000100;
      378: character_line_data <= 'b00001000;
      379: character_line_data <= 'b00010000;
      380: character_line_data <= 'b00100000;
      381: character_line_data <= 'b01000000;
      382: character_line_data <= 'b10000000;
      383: character_line_data <= 'b00000000;
      384: character_line_data <= 'b00111100;
      385: character_line_data <= 'b01000010;
      386: character_line_data <= 'b01000010;
      387: character_line_data <= 'b01000010;
      388: character_line_data <= 'b01000010;
      389: character_line_data <= 'b01000010;
      390: character_line_data <= 'b00111100;
      391: character_line_data <= 'b00000000;
      392: character_line_data <= 'b00010000;
      393: character_line_data <= 'b00110000;
      394: character_line_data <= 'b00010000;
      395: character_line_data <= 'b00010000;
      396: character_line_data <= 'b00010000;
      397: character_line_data <= 'b00010000;
      398: character_line_data <= 'b00111000;
      399: character_line_data <= 'b00000000;
      400: character_line_data <= 'b00111100;
      401: character_line_data <= 'b01000010;
      402: character_line_data <= 'b00000010;
      403: character_line_data <= 'b00001100;
      404: character_line_data <= 'b00110000;
      405: character_line_data <= 'b01000000;
      406: character_line_data <= 'b01111110;
      407: character_line_data <= 'b00000000;
      408: character_line_data <= 'b00111100;
      409: character_line_data <= 'b01000010;
      410: character_line_data <= 'b00000010;
      411: character_line_data <= 'b00011100;
      412: character_line_data <= 'b00000010;
      413: character_line_data <= 'b01000010;
      414: character_line_data <= 'b00111100;
      415: character_line_data <= 'b00000000;
      416: character_line_data <= 'b00000100;
      417: character_line_data <= 'b00001100;
      418: character_line_data <= 'b00010100;
      419: character_line_data <= 'b00100100;
      420: character_line_data <= 'b01000100;
      421: character_line_data <= 'b01111110;
      422: character_line_data <= 'b00000100;
      423: character_line_data <= 'b00000000;
      424: character_line_data <= 'b01111110;
      425: character_line_data <= 'b01000000;
      426: character_line_data <= 'b01111100;
      427: character_line_data <= 'b01000010;
      428: character_line_data <= 'b00000010;
      429: character_line_data <= 'b01000010;
      430: character_line_data <= 'b00111100;
      431: character_line_data <= 'b00000000;
      432: character_line_data <= 'b00111100;
      433: character_line_data <= 'b01000010;
      434: character_line_data <= 'b01000000;
      435: character_line_data <= 'b01111100;
      436: character_line_data <= 'b01000010;
      437: character_line_data <= 'b01000010;
      438: character_line_data <= 'b00111100;
      439: character_line_data <= 'b00000000;
      440: character_line_data <= 'b01111110;
      441: character_line_data <= 'b00000010;
      442: character_line_data <= 'b00000100;
      443: character_line_data <= 'b00001000;
      444: character_line_data <= 'b00001000;
      445: character_line_data <= 'b00010000;
      446: character_line_data <= 'b00010000;
      447: character_line_data <= 'b00000000;
      448: character_line_data <= 'b00111100;
      449: character_line_data <= 'b01000010;
      450: character_line_data <= 'b01000010;
      451: character_line_data <= 'b00111100;
      452: character_line_data <= 'b01000010;
      453: character_line_data <= 'b01000010;
      454: character_line_data <= 'b00111100;
      455: character_line_data <= 'b00000000;
      456: character_line_data <= 'b00111100;
      457: character_line_data <= 'b01000010;
      458: character_line_data <= 'b01000010;
      459: character_line_data <= 'b00111110;
      460: character_line_data <= 'b00000010;
      461: character_line_data <= 'b01000010;
      462: character_line_data <= 'b00111100;
      463: character_line_data <= 'b00000000;
      464: character_line_data <= 'b00000000;
      465: character_line_data <= 'b00110000;
      466: character_line_data <= 'b00110000;
      467: character_line_data <= 'b00000000;
      468: character_line_data <= 'b00110000;
      469: character_line_data <= 'b00110000;
      470: character_line_data <= 'b00000000;
      471: character_line_data <= 'b00000000;
      472: character_line_data <= 'b00000000;
      473: character_line_data <= 'b00110000;
      474: character_line_data <= 'b00110000;
      475: character_line_data <= 'b00000000;
      476: character_line_data <= 'b00110000;
      477: character_line_data <= 'b00010000;
      478: character_line_data <= 'b00100000;
      479: character_line_data <= 'b00000000;
      480: character_line_data <= 'b00000010;
      481: character_line_data <= 'b00000100;
      482: character_line_data <= 'b00001000;
      483: character_line_data <= 'b00010000;
      484: character_line_data <= 'b00001000;
      485: character_line_data <= 'b00000100;
      486: character_line_data <= 'b00000010;
      487: character_line_data <= 'b00000000;
      488: character_line_data <= 'b00000000;
      489: character_line_data <= 'b00000000;
      490: character_line_data <= 'b11111110;
      491: character_line_data <= 'b00000000;
      492: character_line_data <= 'b11111110;
      493: character_line_data <= 'b00000000;
      494: character_line_data <= 'b00000000;
      495: character_line_data <= 'b00000000;
      496: character_line_data <= 'b10000000;
      497: character_line_data <= 'b01000000;
      498: character_line_data <= 'b00100000;
      499: character_line_data <= 'b00010000;
      500: character_line_data <= 'b00100000;
      501: character_line_data <= 'b01000000;
      502: character_line_data <= 'b10000000;
      503: character_line_data <= 'b00000000;
      504: character_line_data <= 'b00111100;
      505: character_line_data <= 'b01000010;
      506: character_line_data <= 'b00000010;
      507: character_line_data <= 'b00001100;
      508: character_line_data <= 'b00010000;
      509: character_line_data <= 'b00000000;
      510: character_line_data <= 'b00010000;
      511: character_line_data <= 'b00000000;
      512: character_line_data <= 'b00111000;
      513: character_line_data <= 'b01000100;
      514: character_line_data <= 'b10011010;
      515: character_line_data <= 'b10101010;
      516: character_line_data <= 'b10110100;
      517: character_line_data <= 'b01000000;
      518: character_line_data <= 'b00111000;
      519: character_line_data <= 'b00000000;
      520: character_line_data <= 'b00010000;
      521: character_line_data <= 'b00101000;
      522: character_line_data <= 'b00101000;
      523: character_line_data <= 'b01000100;
      524: character_line_data <= 'b01111100;
      525: character_line_data <= 'b10000010;
      526: character_line_data <= 'b10000010;
      527: character_line_data <= 'b00000000;
      528: character_line_data <= 'b01111100;
      529: character_line_data <= 'b01000010;
      530: character_line_data <= 'b01000010;
      531: character_line_data <= 'b01111100;
      532: character_line_data <= 'b01000010;
      533: character_line_data <= 'b01000010;
      534: character_line_data <= 'b01111100;
      535: character_line_data <= 'b00000000;
      536: character_line_data <= 'b00011100;
      537: character_line_data <= 'b00100010;
      538: character_line_data <= 'b01000000;
      539: character_line_data <= 'b01000000;
      540: character_line_data <= 'b01000000;
      541: character_line_data <= 'b00100010;
      542: character_line_data <= 'b00011100;
      543: character_line_data <= 'b00000000;
      544: character_line_data <= 'b01111000;
      545: character_line_data <= 'b01000100;
      546: character_line_data <= 'b01000010;
      547: character_line_data <= 'b01000010;
      548: character_line_data <= 'b01000010;
      549: character_line_data <= 'b01000100;
      550: character_line_data <= 'b01111000;
      551: character_line_data <= 'b00000000;
      552: character_line_data <= 'b01111110;
      553: character_line_data <= 'b01000000;
      554: character_line_data <= 'b01000000;
      555: character_line_data <= 'b01111100;
      556: character_line_data <= 'b01000000;
      557: character_line_data <= 'b01000000;
      558: character_line_data <= 'b01111110;
      559: character_line_data <= 'b00000000;
      560: character_line_data <= 'b01111110;
      561: character_line_data <= 'b01000000;
      562: character_line_data <= 'b01000000;
      563: character_line_data <= 'b01111100;
      564: character_line_data <= 'b01000000;
      565: character_line_data <= 'b01000000;
      566: character_line_data <= 'b01000000;
      567: character_line_data <= 'b00000000;
      568: character_line_data <= 'b00011100;
      569: character_line_data <= 'b00100010;
      570: character_line_data <= 'b01000000;
      571: character_line_data <= 'b01001110;
      572: character_line_data <= 'b01000010;
      573: character_line_data <= 'b00100010;
      574: character_line_data <= 'b00011100;
      575: character_line_data <= 'b00000000;
      576: character_line_data <= 'b01000010;
      577: character_line_data <= 'b01000010;
      578: character_line_data <= 'b01000010;
      579: character_line_data <= 'b01111110;
      580: character_line_data <= 'b01000010;
      581: character_line_data <= 'b01000010;
      582: character_line_data <= 'b01000010;
      583: character_line_data <= 'b00000000;
      584: character_line_data <= 'b00111000;
      585: character_line_data <= 'b00010000;
      586: character_line_data <= 'b00010000;
      587: character_line_data <= 'b00010000;
      588: character_line_data <= 'b00010000;
      589: character_line_data <= 'b00010000;
      590: character_line_data <= 'b00111000;
      591: character_line_data <= 'b00000000;
      592: character_line_data <= 'b00000010;
      593: character_line_data <= 'b00000010;
      594: character_line_data <= 'b00000010;
      595: character_line_data <= 'b00000010;
      596: character_line_data <= 'b00000010;
      597: character_line_data <= 'b01000010;
      598: character_line_data <= 'b00111100;
      599: character_line_data <= 'b00000000;
      600: character_line_data <= 'b01000010;
      601: character_line_data <= 'b01000100;
      602: character_line_data <= 'b01001000;
      603: character_line_data <= 'b01010000;
      604: character_line_data <= 'b01101000;
      605: character_line_data <= 'b01000100;
      606: character_line_data <= 'b01000010;
      607: character_line_data <= 'b00000000;
      608: character_line_data <= 'b01000000;
      609: character_line_data <= 'b01000000;
      610: character_line_data <= 'b01000000;
      611: character_line_data <= 'b01000000;
      612: character_line_data <= 'b01000000;
      613: character_line_data <= 'b01000000;
      614: character_line_data <= 'b01111110;
      615: character_line_data <= 'b00000000;
      616: character_line_data <= 'b10000010;
      617: character_line_data <= 'b11000110;
      618: character_line_data <= 'b10101010;
      619: character_line_data <= 'b10101010;
      620: character_line_data <= 'b10010010;
      621: character_line_data <= 'b10010010;
      622: character_line_data <= 'b10000010;
      623: character_line_data <= 'b00000000;
      624: character_line_data <= 'b01000010;
      625: character_line_data <= 'b01100010;
      626: character_line_data <= 'b01010010;
      627: character_line_data <= 'b01001010;
      628: character_line_data <= 'b01000110;
      629: character_line_data <= 'b01000010;
      630: character_line_data <= 'b01000010;
      631: character_line_data <= 'b00000000;
      632: character_line_data <= 'b00011000;
      633: character_line_data <= 'b00100100;
      634: character_line_data <= 'b01000010;
      635: character_line_data <= 'b01000010;
      636: character_line_data <= 'b01000010;
      637: character_line_data <= 'b00100100;
      638: character_line_data <= 'b00011000;
      639: character_line_data <= 'b00000000;
      640: character_line_data <= 'b01111100;
      641: character_line_data <= 'b01000010;
      642: character_line_data <= 'b01000010;
      643: character_line_data <= 'b01111100;
      644: character_line_data <= 'b01000000;
      645: character_line_data <= 'b01000000;
      646: character_line_data <= 'b01000000;
      647: character_line_data <= 'b00000000;
      648: character_line_data <= 'b00011000;
      649: character_line_data <= 'b00100100;
      650: character_line_data <= 'b01000010;
      651: character_line_data <= 'b01000010;
      652: character_line_data <= 'b01001010;
      653: character_line_data <= 'b00100100;
      654: character_line_data <= 'b00011010;
      655: character_line_data <= 'b00000000;
      656: character_line_data <= 'b01111100;
      657: character_line_data <= 'b01000010;
      658: character_line_data <= 'b01000010;
      659: character_line_data <= 'b01111100;
      660: character_line_data <= 'b01001000;
      661: character_line_data <= 'b01000100;
      662: character_line_data <= 'b01000010;
      663: character_line_data <= 'b00000000;
      664: character_line_data <= 'b00111100;
      665: character_line_data <= 'b01000010;
      666: character_line_data <= 'b01000000;
      667: character_line_data <= 'b00111100;
      668: character_line_data <= 'b00000010;
      669: character_line_data <= 'b01000010;
      670: character_line_data <= 'b00111100;
      671: character_line_data <= 'b00000000;
      672: character_line_data <= 'b11111110;
      673: character_line_data <= 'b00010000;
      674: character_line_data <= 'b00010000;
      675: character_line_data <= 'b00010000;
      676: character_line_data <= 'b00010000;
      677: character_line_data <= 'b00010000;
      678: character_line_data <= 'b00010000;
      679: character_line_data <= 'b00000000;
      680: character_line_data <= 'b01000010;
      681: character_line_data <= 'b01000010;
      682: character_line_data <= 'b01000010;
      683: character_line_data <= 'b01000010;
      684: character_line_data <= 'b01000010;
      685: character_line_data <= 'b01000010;
      686: character_line_data <= 'b00111100;
      687: character_line_data <= 'b00000000;
      688: character_line_data <= 'b10000010;
      689: character_line_data <= 'b10000010;
      690: character_line_data <= 'b01000100;
      691: character_line_data <= 'b01000100;
      692: character_line_data <= 'b00101000;
      693: character_line_data <= 'b00101000;
      694: character_line_data <= 'b00010000;
      695: character_line_data <= 'b00000000;
      696: character_line_data <= 'b10000010;
      697: character_line_data <= 'b10010010;
      698: character_line_data <= 'b10010010;
      699: character_line_data <= 'b10101010;
      700: character_line_data <= 'b10101010;
      701: character_line_data <= 'b01000100;
      702: character_line_data <= 'b01000100;
      703: character_line_data <= 'b00000000;
      704: character_line_data <= 'b10000010;
      705: character_line_data <= 'b01000100;
      706: character_line_data <= 'b00101000;
      707: character_line_data <= 'b00010000;
      708: character_line_data <= 'b00101000;
      709: character_line_data <= 'b01000100;
      710: character_line_data <= 'b10000010;
      711: character_line_data <= 'b00000000;
      712: character_line_data <= 'b10000010;
      713: character_line_data <= 'b01000100;
      714: character_line_data <= 'b00101000;
      715: character_line_data <= 'b00010000;
      716: character_line_data <= 'b00010000;
      717: character_line_data <= 'b00010000;
      718: character_line_data <= 'b00010000;
      719: character_line_data <= 'b00000000;
      720: character_line_data <= 'b01111110;
      721: character_line_data <= 'b00000010;
      722: character_line_data <= 'b00000100;
      723: character_line_data <= 'b00001000;
      724: character_line_data <= 'b00010000;
      725: character_line_data <= 'b00100000;
      726: character_line_data <= 'b01111110;
      727: character_line_data <= 'b00000000;
      728: character_line_data <= 'b00001110;
      729: character_line_data <= 'b00001000;
      730: character_line_data <= 'b00001000;
      731: character_line_data <= 'b00001000;
      732: character_line_data <= 'b00001000;
      733: character_line_data <= 'b00001000;
      734: character_line_data <= 'b00001110;
      735: character_line_data <= 'b00000000;
      736: character_line_data <= 'b10000000;
      737: character_line_data <= 'b01000000;
      738: character_line_data <= 'b00100000;
      739: character_line_data <= 'b00010000;
      740: character_line_data <= 'b00001000;
      741: character_line_data <= 'b00000100;
      742: character_line_data <= 'b00000010;
      743: character_line_data <= 'b00000000;
      744: character_line_data <= 'b11100000;
      745: character_line_data <= 'b00100000;
      746: character_line_data <= 'b00100000;
      747: character_line_data <= 'b00100000;
      748: character_line_data <= 'b00100000;
      749: character_line_data <= 'b00100000;
      750: character_line_data <= 'b11100000;
      751: character_line_data <= 'b00000000;
      752: character_line_data <= 'b00010000;
      753: character_line_data <= 'b00101000;
      754: character_line_data <= 'b01000100;
      755: character_line_data <= 'b00000000;
      756: character_line_data <= 'b00000000;
      757: character_line_data <= 'b00000000;
      758: character_line_data <= 'b00000000;
      759: character_line_data <= 'b00000000;
      760: character_line_data <= 'b00000000;
      761: character_line_data <= 'b00000000;
      762: character_line_data <= 'b00000000;
      763: character_line_data <= 'b00000000;
      764: character_line_data <= 'b00000000;
      765: character_line_data <= 'b00000000;
      766: character_line_data <= 'b11111110;
      767: character_line_data <= 'b00000000;
      768: character_line_data <= 'b10000000;
      769: character_line_data <= 'b01000000;
      770: character_line_data <= 'b00100000;
      771: character_line_data <= 'b00000000;
      772: character_line_data <= 'b00000000;
      773: character_line_data <= 'b00000000;
      774: character_line_data <= 'b00000000;
      775: character_line_data <= 'b00000000;
      776: character_line_data <= 'b00000000;
      777: character_line_data <= 'b00000000;
      778: character_line_data <= 'b00111000;
      779: character_line_data <= 'b00000100;
      780: character_line_data <= 'b00111100;
      781: character_line_data <= 'b01000100;
      782: character_line_data <= 'b00111100;
      783: character_line_data <= 'b00000000;
      784: character_line_data <= 'b01000000;
      785: character_line_data <= 'b01000000;
      786: character_line_data <= 'b01011000;
      787: character_line_data <= 'b01100100;
      788: character_line_data <= 'b01000100;
      789: character_line_data <= 'b01000100;
      790: character_line_data <= 'b01111000;
      791: character_line_data <= 'b00000000;
      792: character_line_data <= 'b00000000;
      793: character_line_data <= 'b00000000;
      794: character_line_data <= 'b00111000;
      795: character_line_data <= 'b01000100;
      796: character_line_data <= 'b01000000;
      797: character_line_data <= 'b01000100;
      798: character_line_data <= 'b00111000;
      799: character_line_data <= 'b00000000;
      800: character_line_data <= 'b00000100;
      801: character_line_data <= 'b00000100;
      802: character_line_data <= 'b00110100;
      803: character_line_data <= 'b01001100;
      804: character_line_data <= 'b01000100;
      805: character_line_data <= 'b01000100;
      806: character_line_data <= 'b00111100;
      807: character_line_data <= 'b00000000;
      808: character_line_data <= 'b00000000;
      809: character_line_data <= 'b00000000;
      810: character_line_data <= 'b00111000;
      811: character_line_data <= 'b01000100;
      812: character_line_data <= 'b01111100;
      813: character_line_data <= 'b01000000;
      814: character_line_data <= 'b00111000;
      815: character_line_data <= 'b00000000;
      816: character_line_data <= 'b00001100;
      817: character_line_data <= 'b00010000;
      818: character_line_data <= 'b00111000;
      819: character_line_data <= 'b00010000;
      820: character_line_data <= 'b00010000;
      821: character_line_data <= 'b00010000;
      822: character_line_data <= 'b00010000;
      823: character_line_data <= 'b00000000;
      824: character_line_data <= 'b00000000;
      825: character_line_data <= 'b00000000;
      826: character_line_data <= 'b00111100;
      827: character_line_data <= 'b01000100;
      828: character_line_data <= 'b00111100;
      829: character_line_data <= 'b00000100;
      830: character_line_data <= 'b00111000;
      831: character_line_data <= 'b00000000;
      832: character_line_data <= 'b01000000;
      833: character_line_data <= 'b01000000;
      834: character_line_data <= 'b01011000;
      835: character_line_data <= 'b01100100;
      836: character_line_data <= 'b01000100;
      837: character_line_data <= 'b01000100;
      838: character_line_data <= 'b01000100;
      839: character_line_data <= 'b00000000;
      840: character_line_data <= 'b00010000;
      841: character_line_data <= 'b00000000;
      842: character_line_data <= 'b00010000;
      843: character_line_data <= 'b00010000;
      844: character_line_data <= 'b00010000;
      845: character_line_data <= 'b00010000;
      846: character_line_data <= 'b00010000;
      847: character_line_data <= 'b00000000;
      848: character_line_data <= 'b00001000;
      849: character_line_data <= 'b00000000;
      850: character_line_data <= 'b00001000;
      851: character_line_data <= 'b00001000;
      852: character_line_data <= 'b00001000;
      853: character_line_data <= 'b01001000;
      854: character_line_data <= 'b00110000;
      855: character_line_data <= 'b00000000;
      856: character_line_data <= 'b00100000;
      857: character_line_data <= 'b00100000;
      858: character_line_data <= 'b00100100;
      859: character_line_data <= 'b00101000;
      860: character_line_data <= 'b00110000;
      861: character_line_data <= 'b00101000;
      862: character_line_data <= 'b00100100;
      863: character_line_data <= 'b00000000;
      864: character_line_data <= 'b00110000;
      865: character_line_data <= 'b00010000;
      866: character_line_data <= 'b00010000;
      867: character_line_data <= 'b00010000;
      868: character_line_data <= 'b00010000;
      869: character_line_data <= 'b00010000;
      870: character_line_data <= 'b00010000;
      871: character_line_data <= 'b00000000;
      872: character_line_data <= 'b00000000;
      873: character_line_data <= 'b00000000;
      874: character_line_data <= 'b01101000;
      875: character_line_data <= 'b01010100;
      876: character_line_data <= 'b01010100;
      877: character_line_data <= 'b01010100;
      878: character_line_data <= 'b01010100;
      879: character_line_data <= 'b00000000;
      880: character_line_data <= 'b00000000;
      881: character_line_data <= 'b00000000;
      882: character_line_data <= 'b01011000;
      883: character_line_data <= 'b01100100;
      884: character_line_data <= 'b01000100;
      885: character_line_data <= 'b01000100;
      886: character_line_data <= 'b01000100;
      887: character_line_data <= 'b00000000;
      888: character_line_data <= 'b00000000;
      889: character_line_data <= 'b00000000;
      890: character_line_data <= 'b00111000;
      891: character_line_data <= 'b01000100;
      892: character_line_data <= 'b01000100;
      893: character_line_data <= 'b01000100;
      894: character_line_data <= 'b00111000;
      895: character_line_data <= 'b00000000;
      896: character_line_data <= 'b00000000;
      897: character_line_data <= 'b00000000;
      898: character_line_data <= 'b01111000;
      899: character_line_data <= 'b01000100;
      900: character_line_data <= 'b01111000;
      901: character_line_data <= 'b01000000;
      902: character_line_data <= 'b01000000;
      903: character_line_data <= 'b00000000;
      904: character_line_data <= 'b00000000;
      905: character_line_data <= 'b00000000;
      906: character_line_data <= 'b00111100;
      907: character_line_data <= 'b01000100;
      908: character_line_data <= 'b00111100;
      909: character_line_data <= 'b00000100;
      910: character_line_data <= 'b00000100;
      911: character_line_data <= 'b00000000;
      912: character_line_data <= 'b00000000;
      913: character_line_data <= 'b00000000;
      914: character_line_data <= 'b01011000;
      915: character_line_data <= 'b01100100;
      916: character_line_data <= 'b01000000;
      917: character_line_data <= 'b01000000;
      918: character_line_data <= 'b01000000;
      919: character_line_data <= 'b00000000;
      920: character_line_data <= 'b00000000;
      921: character_line_data <= 'b00000000;
      922: character_line_data <= 'b00111100;
      923: character_line_data <= 'b01000000;
      924: character_line_data <= 'b00111000;
      925: character_line_data <= 'b00000100;
      926: character_line_data <= 'b01111000;
      927: character_line_data <= 'b00000000;
      928: character_line_data <= 'b00000000;
      929: character_line_data <= 'b00100000;
      930: character_line_data <= 'b01111000;
      931: character_line_data <= 'b00100000;
      932: character_line_data <= 'b00100000;
      933: character_line_data <= 'b00100100;
      934: character_line_data <= 'b00011000;
      935: character_line_data <= 'b00000000;
      936: character_line_data <= 'b00000000;
      937: character_line_data <= 'b00000000;
      938: character_line_data <= 'b01000100;
      939: character_line_data <= 'b01000100;
      940: character_line_data <= 'b01000100;
      941: character_line_data <= 'b01001100;
      942: character_line_data <= 'b00110100;
      943: character_line_data <= 'b00000000;
      944: character_line_data <= 'b00000000;
      945: character_line_data <= 'b00000000;
      946: character_line_data <= 'b01000100;
      947: character_line_data <= 'b01000100;
      948: character_line_data <= 'b00101000;
      949: character_line_data <= 'b00101000;
      950: character_line_data <= 'b00010000;
      951: character_line_data <= 'b00000000;
      952: character_line_data <= 'b00000000;
      953: character_line_data <= 'b00000000;
      954: character_line_data <= 'b01000100;
      955: character_line_data <= 'b01010100;
      956: character_line_data <= 'b01010100;
      957: character_line_data <= 'b00101000;
      958: character_line_data <= 'b00101000;
      959: character_line_data <= 'b00000000;
      960: character_line_data <= 'b00000000;
      961: character_line_data <= 'b00000000;
      962: character_line_data <= 'b01000100;
      963: character_line_data <= 'b00101000;
      964: character_line_data <= 'b00010000;
      965: character_line_data <= 'b00101000;
      966: character_line_data <= 'b01000100;
      967: character_line_data <= 'b00000000;
      968: character_line_data <= 'b00000000;
      969: character_line_data <= 'b00000000;
      970: character_line_data <= 'b01000100;
      971: character_line_data <= 'b00101000;
      972: character_line_data <= 'b00101000;
      973: character_line_data <= 'b00010000;
      974: character_line_data <= 'b01100000;
      975: character_line_data <= 'b00000000;
      976: character_line_data <= 'b00000000;
      977: character_line_data <= 'b00000000;
      978: character_line_data <= 'b01111100;
      979: character_line_data <= 'b00001000;
      980: character_line_data <= 'b00010000;
      981: character_line_data <= 'b00100000;
      982: character_line_data <= 'b01111100;
      983: character_line_data <= 'b00000000;
      984: character_line_data <= 'b00000110;
      985: character_line_data <= 'b00001000;
      986: character_line_data <= 'b00001000;
      987: character_line_data <= 'b00010000;
      988: character_line_data <= 'b00001000;
      989: character_line_data <= 'b00001000;
      990: character_line_data <= 'b00000110;
      991: character_line_data <= 'b00000000;
      992: character_line_data <= 'b00010000;
      993: character_line_data <= 'b00010000;
      994: character_line_data <= 'b00010000;
      995: character_line_data <= 'b00010000;
      996: character_line_data <= 'b00010000;
      997: character_line_data <= 'b00010000;
      998: character_line_data <= 'b00010000;
      999: character_line_data <= 'b00000000;
      1000: character_line_data <= 'b11000000;
      1001: character_line_data <= 'b00100000;
      1002: character_line_data <= 'b00100000;
      1003: character_line_data <= 'b00010000;
      1004: character_line_data <= 'b00100000;
      1005: character_line_data <= 'b00100000;
      1006: character_line_data <= 'b11000000;
      1007: character_line_data <= 'b00000000;
      1008: character_line_data <= 'b00000000;
      1009: character_line_data <= 'b00000000;
      1010: character_line_data <= 'b01100000;
      1011: character_line_data <= 'b10010010;
      1012: character_line_data <= 'b00001100;
      1013: character_line_data <= 'b00000000;
      1014: character_line_data <= 'b00000000;
      1015: character_line_data <= 'b00000000;
      1016: character_line_data <= 'b00000000;
      1017: character_line_data <= 'b00000000;
      1018: character_line_data <= 'b00000000;
      1019: character_line_data <= 'b00000000;
      1020: character_line_data <= 'b00000000;
      1021: character_line_data <= 'b00000000;
      1022: character_line_data <= 'b00000000;
      1023: character_line_data <= 'b00000000;
    endcase
  end
endmodule

`timescale 1ns / 1ps

module index();
endmodule

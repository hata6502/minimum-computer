module index();
endmodule
